StartDeckInitial
1
JS
2
KC
3
5C
4
2H
5
9S
6
AS
7
3H
8
6C
9
8D
10
AC
11
10S
12
5H
13
2D
14
KD
15
7D
16
8C
17
3S
18
AD
19
7S
20
5S
21
QD
22
AH
23
8S
24
3D
25
7H
26
QH
27
5D
28
7C
29
4H
30
KH
31
4D
32
10D
33
JC
34
JH
35
10C
36
JD
37
4S
38
10H
39
6H
40
3C
41
2S
42
9H
43
KS
44
6S
45
4C
46
8H
47
9C
48
QS
49
6D
50
QC
51
2C
52
9D
StartDeck
49
6D
44
6S
33
JC
28
7C
17
3S
38
10H
1
JS
22
AH
11
10S
6
AS
46
8H
41
2S
30
KH
51
2C
14
KD
35
10C
24
3D
19
7S
8
6C
3
5C
43
KS
13
2D
27
5D
48
QS
37
4S
32
10D
21
QD
16
8C
5
9S
26
QH
40
3C
10
AC
50
QC
45
4C
34
JH
29
4H
18
AD
39
6H
2
KC
23
8S
12
5H
7
3H
47
9C
42
9H
31
4D
52
9D
15
7D
36
JD
25
7H
20
5S
9
8D
4
2H
TargetDeck
49
6D
44
6S
33
JC
28
7C
17
3S
38
10H
1
JS
22
AH
11
10S
6
AS
46
8H
41
2S
30
KH
51
2C
14
KD
35
10C
24
3D
19
7S
8
6C
3
5C
43
KS
13
2D
27
5D
48
QS
37
4S
32
10D
21
QD
16
8C
5
9S
26
QH
40
3C
10
AC
50
QC
45
4C
34
JH
29
4H
18
AD
39
6H
2
KC
23
8S
12
5H
7
3H
47
9C
42
9H
31
4D
52
9D
15
7D
36
JD
25
7H
20
5S
9
8D
4
2H
StartDeckName
Aronson.svf
TargetDeckName
AronsonChanged3.svf
SearchLevels
5
CutDeckPrecise
8
45
52
1
0
RunSingleCards
0
0
0
0
0
RunSingleCardsInv
0
0
0
0
0
SearchMoveCard
0
0
0
0
0
0
0
SearchShiftTopBlock
0
0
0
0
0
0
0
SearchShiftTopBlockInv
0
0
0
0
0
0
0
SearchOutFaro
1
SearchOutFaroInverse
0
SearchOutFaroSpecialTop
0
0
0
0
0
0
0
SearchOutFaroSpecialTopInv
0
0
0
0
0
0
0
SearchOutFaroSpecialBottom
0
0
0
0
0
0
0
SearchOutFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchInFaro
1
SearchInFaroInverse
0
SearchInFaroSpecialTop
0
0
0
0
0
0
0
SearchInFaroSpecialTopInv
0
0
0
0
0
0
0
SearchInFaroSpecialBottom
0
0
0
0
0
0
0
SearchInFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchLevelCounter(x)
9
9
10
10
9
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
MatchFound
1
NoMatchFound
0
SearchStartDeckSet
1
SearchTargetDeckSet
1
SearchCurrentLevel
5
SearchCurrentLevelRestart
0
SearchProcessing
False
SearchProgressCounter
332
SearchElapsedTime
23.765625
SearchSpecialName
CutDeckPrecise
SearchSessionTransferred
0
SearchingMode
False
SearchCounter
11
SearchContinueReady
0
SearchCounterMax
10
SearchParseError
False
SearchMatchStartCard
1
SearchMatchEndCard
52
WholeDeckMatch
True
PartialDeckMatch
False
ThresholdMatchCards
0
TrapThreshold
False
WholeDeckMatchSet
True
PartialMatchFound
0
ContinueSearchToggle(0)
False
ContinueSearchToggle(1)
False
TimerResult
23 secs
ProgressLabel

SearchTimeLabel
21 secs 
ManipulationsLabel
10
TrapFileWhole

TrapFileWholeFinal

TrapFileFinal

TrapPathWhole

TrapPathWholeFinal

TrapPathFinal

TrapFilePartial

TrapFilePartialFinal

TrapPathPartial

TrapPathPartialFinal

SuspendTrapWhole

SuspendTrapPartial

SuspendTrapWholeFinal

SuspendTrapPartialFinal

SuspendTrapFinal
True
PartialDeckMatchStart

PartialDeckMatchEnd

PartialDeckMatchThresholdCards

PartialDeckMatchThresholdCheck
0
WholeDeckMatchThresholdCards
0
WholeDeckMatchThresholdCheck
0
SolutionResults
OutFaro
OutFaro
InFaro
InFaro
OutFaro
