StartDeckInitial
1
JS
2
KC
3
5C
4
2H
5
9S
6
AS
7
3H
8
6C
9
8D
10
AC
11
10S
12
5H
13
2D
14
KD
15
7D
16
8C
17
3S
18
AD
19
7S
20
5S
21
QD
22
AH
23
8S
24
3D
25
7H
26
QH
27
5D
28
7C
29
4H
30
KH
31
4D
32
10D
33
JC
34
JH
35
10C
36
JD
37
4S
38
10H
39
6H
40
3C
41
2S
42
9H
43
KS
44
6S
45
4C
46
8H
47
9C
48
QS
49
6D
50
QC
51
2C
52
9D
StartDeck
27
5D
1
JS
28
7C
2
KC
29
4H
3
5C
30
KH
4
2H
31
4D
5
9S
32
10D
6
AS
33
JC
7
3H
34
JH
8
6C
35
10C
9
8D
36
JD
10
AC
37
4S
11
10S
38
10H
12
5H
39
6H
13
2D
40
3C
14
KD
41
2S
15
7D
42
9H
16
8C
43
KS
17
3S
44
6S
18
AD
45
4C
19
7S
46
8H
20
5S
47
9C
21
QD
48
QS
22
AH
49
6D
23
8S
50
QC
24
3D
51
2C
25
7H
52
9D
26
QH
TargetDeck
15
7D
34
JH
36
JD
31
4D
21
QD
28
7C
40
3C
46
8H
23
8S
8
6C
30
KH
7
3H
52
9D
22
AH
39
6H
24
3D
27
5D
44
6S
50
QC
49
6D
45
4C
47
9C
10
AC
35
10C
9
8D
25
7H
32
10D
19
7S
6
AS
33
JC
41
2S
37
4S
5
9S
1
JS
14
KD
16
8C
29
4H
17
3S
42
9H
11
10S
13
2D
2
KC
51
2C
18
AD
3
5C
4
2H
20
5S
26
QH
43
KS
12
5H
48
QS
38
10H
StartDeckName
Aronson.svf
TargetDeckName
AronsonChanged4.svf
SearchLevels
5
CutDeckPrecise
8
45
52
1
0
RunSingleCards
0
0
0
0
0
RunSingleCardsInv
0
0
0
0
0
SearchMoveCard
0
0
0
0
0
0
0
SearchShiftTopBlock
0
0
0
0
0
0
0
SearchShiftTopBlockInv
0
0
0
0
0
0
0
SearchOutFaro
1
SearchOutFaroInverse
0
SearchOutFaroSpecialTop
0
0
0
0
0
0
0
SearchOutFaroSpecialTopInv
0
0
0
0
0
0
0
SearchOutFaroSpecialBottom
0
0
0
0
0
0
0
SearchOutFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchInFaro
1
SearchInFaroInverse
0
SearchInFaroSpecialTop
0
0
0
0
0
0
0
SearchInFaroSpecialTopInv
0
0
0
0
0
0
0
SearchInFaroSpecialBottom
0
0
0
0
0
0
0
SearchInFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchLevelCounter(x)
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
MatchFound
0
NoMatchFound
1
SearchStartDeckSet
1
SearchTargetDeckSet
1
SearchCurrentLevel
6
SearchCurrentLevelRestart
0
SearchProcessing
False
SearchProgressCounter
340
SearchElapsedTime
21.078125
SearchSpecialName
CutDeckPrecise
SearchSessionTransferred
0
SearchingMode
False
SearchCounter
11
SearchContinueReady
0
SearchCounterMax
10
SearchParseError
False
SearchMatchStartCard
1
SearchMatchEndCard
52
WholeDeckMatch
True
PartialDeckMatch
False
ThresholdMatchCards
0
TrapThreshold
False
WholeDeckMatchSet
True
PartialMatchFound
0
ContinueSearchToggle(0)
False
ContinueSearchToggle(1)
False
TimerResult
21 secs
ProgressLabel

SearchTimeLabel
21 secs 
ManipulationsLabel
10
TrapFileWhole

TrapFileWholeFinal

TrapFileFinal

TrapPathWhole

TrapPathWholeFinal

TrapPathFinal

TrapFilePartial

TrapFilePartialFinal

TrapPathPartial

TrapPathPartialFinal

SuspendTrapWhole

SuspendTrapPartial

SuspendTrapWholeFinal

SuspendTrapPartialFinal

SuspendTrapFinal
True
PartialDeckMatchStart

PartialDeckMatchEnd

PartialDeckMatchThresholdCards

PartialDeckMatchThresholdCheck
0
WholeDeckMatchThresholdCards
0
WholeDeckMatchThresholdCheck
0
