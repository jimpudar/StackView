StartDeckInitial
1
JS
2
KC
3
5C
4
2H
5
9S
6
AS
7
3H
8
6C
9
8D
10
AC
11
10S
12
5H
13
2D
14
KD
15
7D
16
8C
17
3S
18
AD
19
7S
20
5S
21
QD
22
AH
23
8S
24
3D
25
7H
26
QH
27
5D
28
7C
29
4H
30
KH
31
4D
32
10D
33
JC
34
JH
35
10C
36
JD
37
4S
38
10H
39
6H
40
3C
41
2S
42
9H
43
KS
44
6S
45
4C
46
8H
47
9C
48
QS
49
6D
50
QC
51
2C
52
9D
StartDeck








































































































TargetDeck
13
2D
9
8D
5
9S
1
JS
29
4H
25
7H
21
QD
17
3S
45
4C
41
2S
37
4S
33
JC
10
AC
6
AS
2
KC
49
6D
26
QH
22
AH
18
AD
14
KD
42
9H
38
10H
34
JH
30
KH
7
3H
3
5C
50
QC
46
8H
23
8S
19
7S
15
7D
11
10S
39
6H
35
10C
31
4D
27
5D
4
2H
51
2C
47
9C
43
KS
20
5S
16
8C
12
5H
8
6C
36
JD
32
10D
28
7C
24
3D
52
9D
48
QS
44
6S
40
3C
StartDeckName
Aronson.svf
TargetDeckName
AronsonChanged.svf
SearchLevels
5
CutDeckPrecise
5
48
52
1
0
RunSingleCards
0
0
0
0
0
RunSingleCardsInv
0
0
0
0
0
SearchMoveCard
0
0
0
0
0
0
0
SearchShiftTopBlock
0
0
0
0
0
0
0
SearchShiftTopBlockInv
0
0
0
0
0
0
0
SearchOutFaro
1
SearchOutFaroInverse
0
SearchOutFaroSpecialTop
0
0
0
0
0
0
0
SearchOutFaroSpecialTopInv
0
0
0
0
0
0
0
SearchOutFaroSpecialBottom
0
0
0
0
0
0
0
SearchOutFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchInFaro
1
SearchInFaroInverse
0
SearchInFaroSpecialTop
0
0
0
0
0
0
0
SearchInFaroSpecialTopInv
0
0
0
0
0
0
0
SearchInFaroSpecialBottom
0
0
0
0
0
0
0
SearchInFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchLevelCounter(x)
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
0
MatchFound
0
SearchStartDeckSet
1
SearchTargetDeckSet
1
SearchCurrentLevel
0
SearchCurrentLevelRestart
0
SearchProcessing
False
SearchProgressCounter
0
SearchElapsedTime
0
SearchSpecialName
CutDeckPrecise
SearchSessionTransferred
0
SearchingMode
False
SearchCounter
1
SearchContinueReady
0
SearchCounterMax
7
SearchParseError
False
SearchMatchStartCard
1
SearchMatchEndCard
52
WholeDeckMatch
True
PartialDeckMatch
False
ThresholdMatchCards
0
TrapThreshold
False
WholeDeckMatchSet
True
PartialMatchFound
0
ContinueSearchToggle(0)
False
ContinueSearchToggle(1)
False
TimerResult

ProgressLabel

SearchTimeLabel
4 secs 
ManipulationsLabel
7
TrapFileWhole

TrapFileWholeFinal

TrapFileFinal

TrapPathWhole

TrapPathWholeFinal

TrapPathFinal

TrapFilePartial

TrapFilePartialFinal

TrapPathPartial

TrapPathPartialFinal

SuspendTrapWhole

SuspendTrapPartial

SuspendTrapWholeFinal

SuspendTrapPartialFinal

SuspendTrapFinal
True
PartialDeckMatchStart

PartialDeckMatchEnd

PartialDeckMatchThresholdCards

PartialDeckMatchThresholdCheck
0
WholeDeckMatchThresholdCards
0
WholeDeckMatchThresholdCheck
0
