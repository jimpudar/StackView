StartDeckInitial
1
JS
2
KC
3
5C
4
2H
5
9S
6
AS
7
3H
8
6C
9
8D
10
AC
11
10S
12
5H
13
2D
14
KD
15
7D
16
8C
17
3S
18
AD
19
7S
20
5S
21
QD
22
AH
23
8S
24
3D
25
7H
26
QH
27
5D
28
7C
29
4H
30
KH
31
4D
32
10D
33
JC
34
JH
35
10C
36
JD
37
4S
38
10H
39
6H
40
3C
41
2S
42
9H
43
KS
44
6S
45
4C
46
8H
47
9C
48
QS
49
6D
50
QC
51
2C
52
9D
StartDeck
48
QS
23
8S
41
2S
16
8C
34
JH
1
JS
27
5D
7
3H
25
7H
51
2C
18
AD
44
6S
11
10S
29
4H
4
2H
22
AH
40
3C
15
7D
33
JC
8
6C
39
6H
6
AS
32
10D
50
QC
17
3S
43
KS
10
AC
36
JD
3
5C
21
QD
47
9C
14
KD
45
4C
20
5S
38
10H
13
2D
31
4D
49
6D
24
3D
42
9H
9
8D
35
10C
2
KC
28
7C
46
8H
26
QH
52
9D
19
7S
37
4S
12
5H
30
KH
5
9S
TargetDeck
48
QS
23
8S
41
2S
16
8C
34
JH
1
JS
27
5D
7
3H
25
7H
51
2C
18
AD
44
6S
11
10S
29
4H
4
2H
22
AH
40
3C
15
7D
33
JC
8
6C
39
6H
6
AS
32
10D
50
QC
17
3S
43
KS
10
AC
36
JD
3
5C
21
QD
47
9C
14
KD
45
4C
20
5S
38
10H
13
2D
31
4D
49
6D
24
3D
42
9H
9
8D
35
10C
2
KC
28
7C
46
8H
26
QH
52
9D
19
7S
37
4S
12
5H
30
KH
5
9S
StartDeckName
Aronson.svf
TargetDeckName
AronsonChanged2.svf
SearchLevels
9
CutDeckPrecise
2
51
52
1
0
RunSingleCards
0
0
0
0
0
RunSingleCardsInv
0
0
0
0
0
SearchMoveCard
0
0
0
0
0
0
0
SearchShiftTopBlock
0
0
0
0
0
0
0
SearchShiftTopBlockInv
0
0
0
0
0
0
0
SearchOutFaro
1
SearchOutFaroInverse
0
SearchOutFaroSpecialTop
0
0
0
0
0
0
0
SearchOutFaroSpecialTopInv
0
0
0
0
0
0
0
SearchOutFaroSpecialBottom
0
0
0
0
0
0
0
SearchOutFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchInFaro
1
SearchInFaroInverse
0
SearchInFaroSpecialTop
0
0
0
0
0
0
0
SearchInFaroSpecialTopInv
0
0
0
0
0
0
0
SearchInFaroSpecialBottom
0
0
0
0
0
0
0
SearchInFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchLevelCounter(x)
3
3
3
4
4
4
3
3
3
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
MatchFound
1
SearchStartDeckSet
1
SearchTargetDeckSet
1
SearchCurrentLevel
9
SearchCurrentLevelRestart
5
SearchProcessing
False
SearchProgressCounter
34
SearchElapsedTime
62.84375
SearchSpecialName
CutDeckPrecise
SearchSessionTransferred
0
SearchingMode
False
SearchCounter
5
SearchContinueReady
0
SearchCounterMax
4
SearchParseError
False
SearchMatchStartCard
1
SearchMatchEndCard
52
WholeDeckMatch
True
PartialDeckMatch
False
ThresholdMatchCards
0
TrapThreshold
False
WholeDeckMatchSet
True
PartialMatchFound
0
ContinueSearchToggle(0)
False
ContinueSearchToggle(1)
False
TimerResult
1 min 2 secs
ProgressLabel

SearchTimeLabel
1 min 20 secs 
ManipulationsLabel
4
TrapFileWhole

TrapFileWholeFinal

TrapFileFinal

TrapPathWhole

TrapPathWholeFinal

TrapPathFinal

TrapFilePartial

TrapFilePartialFinal

TrapPathPartial

TrapPathPartialFinal

SuspendTrapWhole

SuspendTrapPartial

SuspendTrapWholeFinal

SuspendTrapPartialFinal

SuspendTrapFinal
True
PartialDeckMatchStart

PartialDeckMatchEnd

PartialDeckMatchThresholdCards

PartialDeckMatchThresholdCheck
0
WholeDeckMatchThresholdCards
0
WholeDeckMatchThresholdCheck
0
