StartDeckInitial
1
JS
2
KC
3
5C
4
2H
5
9S
6
AS
7
3H
8
6C
9
8D
10
AC
11
10S
12
5H
13
2D
14
KD
15
7D
16
8C
17
3S
18
AD
19
7S
20
5S
21
QD
22
AH
23
8S
24
3D
25
7H
26
QH
27
5D
28
7C
29
4H
30
KH
31
4D
32
10D
33
JC
34
JH
35
10C
36
JD
37
4S
38
10H
39
6H
40
3C
41
2S
42
9H
43
KS
44
6S
45
4C
46
8H
47
9C
48
QS
49
6D
50
QC
51
2C
52
9D
StartDeck
38
10H
39
6H
40
3C
41
2S
42
9H
43
KS
44
6S
45
4C
46
8H
47
9C
48
QS
49
6D
50
QC
51
2C
52
9D
1
JS
2
KC
3
5C
4
2H
5
9S
6
AS
7
3H
8
6C
9
8D
10
AC
11
10S
12
5H
13
2D
14
KD
15
7D
16
8C
17
3S
18
AD
19
7S
20
5S
21
QD
22
AH
23
8S
24
3D
25
7H
26
QH
27
5D
28
7C
29
4H
30
KH
31
4D
32
10D
33
JC
34
JH
35
10C
36
JD
37
4S
TargetDeck
11
10S
43
KS
24
3D
4
2H
37
4S
50
QC
45
4C
36
JD
12
5H
26
QH
47
9C
25
7H
32
10D
5
9S
33
JC
49
6D
17
3S
15
7D
35
10C
2
KC
18
AD
34
JH
10
AC
48
QS
41
2S
51
2C
39
6H
52
9D
23
8S
27
5D
20
5S
30
KH
6
AS
13
2D
44
6S
21
QD
22
AH
7
3H
9
8D
8
6C
40
3C
16
8C
31
4D
46
8H
14
KD
19
7S
1
JS
38
10H
29
4H
42
9H
3
5C
28
7C
StartDeckName
Aronson.svf
TargetDeckName
AronsonChanged2.svf
SearchLevels
5
CutDeckPrecise
13
40
52
1
0
RunSingleCards
0
0
0
0
0
RunSingleCardsInv
0
0
0
0
0
SearchMoveCard
0
0
0
0
0
0
0
SearchShiftTopBlock
0
0
0
0
0
0
0
SearchShiftTopBlockInv
0
0
0
0
0
0
0
SearchOutFaro
1
SearchOutFaroInverse
0
SearchOutFaroSpecialTop
0
0
0
0
0
0
0
SearchOutFaroSpecialTopInv
0
0
0
0
0
0
0
SearchOutFaroSpecialBottom
0
0
0
0
0
0
0
SearchOutFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchInFaro
0
SearchInFaroInverse
0
SearchInFaroSpecialTop
0
0
0
0
0
0
0
SearchInFaroSpecialTopInv
0
0
0
0
0
0
0
SearchInFaroSpecialBottom
0
0
0
0
0
0
0
SearchInFaroSpecialBottomInv
0
0
0
0
0
0
0
SearchLevelCounter(x)
1
12
11
2
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
MatchFound
0
SearchStartDeckSet
1
SearchTargetDeckSet
1
SearchCurrentLevel
4
SearchCurrentLevelRestart
4
SearchProcessing
False
SearchProgressCounter
0
SearchElapsedTime
0.9375
SearchSpecialName
CutDeckPrecise
SearchSessionTransferred
0
SearchingMode
False
SearchCounter
15
SearchContinueReady
1
SearchCounterMax
14
SearchParseError
False
SearchMatchStartCard
1
SearchMatchEndCard
10
WholeDeckMatch
False
PartialDeckMatch
True
ThresholdMatchCards
5
TrapThreshold
True
WholeDeckMatchSet
False
PartialMatchFound
0
ContinueSearchToggle(0)
True
ContinueSearchToggle(1)
False
TimerResult
0 secs
ProgressLabel
4 [1,12,11,2]
SearchTimeLabel
2 mins 24 secs 
ManipulationsLabel
14
TrapFileWhole

TrapFileWholeFinal

TrapFileFinal

TrapPathWhole

TrapPathWholeFinal

TrapPathFinal

TrapFilePartial

TrapFilePartialFinal

TrapPathPartial

TrapPathPartialFinal

SuspendTrapWhole

SuspendTrapPartial
True
SuspendTrapWholeFinal

SuspendTrapPartialFinal
True
SuspendTrapFinal
True
PartialDeckMatchStart
1
PartialDeckMatchEnd
10
PartialDeckMatchThresholdCards
5
PartialDeckMatchThresholdCheck
1
WholeDeckMatchThresholdCards

WholeDeckMatchThresholdCheck
0
